module and2_primitive (x, y, f);
	input x, y;
	output f;
	
	and INS0 (f, x, y);
endmodule
